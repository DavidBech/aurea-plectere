
module top_test;

logic clk;
logic reset_n;

aurea_plectere #(

) u_dut (
    .clk    (clk    ),
    .reset_n(reset_n)
);






endmodule

