
module aurea_plectere #(


) (
    input logic clk,
    input logic reset_n

);

endmodule

